// CODEC Environment

`include "clock_and_reset_bfm_env.sv"
`include "i2s_bfm_env.sv"
`include "axi4_lite_bfm_env.sv"
`include "codec_unit_top_pkg.svh"