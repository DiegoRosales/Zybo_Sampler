
// TODO Automate this
package codec_unit_top_reg_model_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "codec_registers_uvm_reg_model.sv"
endpackage