// clock_and_reset Verification IP

`include "clock_and_reset_if.svh"
`include "clock_and_reset_bfm_pkg.svh"