// All the testcases

`include "codec_unit_top_base_test.sv"
`include "codec_unit_top_testcase_1.sv"