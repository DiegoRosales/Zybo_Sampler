// Testbench package

package codec_unit_top_pkg;
  // Mandatory UVM
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import i2s_bfm_pkg::*;

  `include "codec_unit_top_base_test_env.svh"
  `include "codec_registers_uvm_reg_model.sv"

endpackage