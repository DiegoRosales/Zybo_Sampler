// I2S Verification IP

`include "i2s_if.svh"
`include "i2s_bfm_pkg.svh"