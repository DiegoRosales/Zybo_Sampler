// clock_and_reset Interface definition for Verification

interface clock_and_reset_if;

  bit clock;
  bit reset;

endinterface //clock_and_reset_if