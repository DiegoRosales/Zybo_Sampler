// CODEC Environment

`include "codec_unit_top_pkg.svh"