// Testbench package

package codec_unit_top_pkg;
  import uvm_pkg::*;


endpackage