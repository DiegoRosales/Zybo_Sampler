/////////////////////////////////////
// AXI4-Lite BFM Environment
/////////////////////////////////////

`include "axi4_lite_if.sv"
`include "axi4_lite_bfm_pkg.sv"